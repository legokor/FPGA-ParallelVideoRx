`timescale 1ns / 1ps

module ov5642_interface(
    input pclk,
    input xclk,
    input href,
    input vsync,
    input [9:0] data,
    output pwdn
    );
    
    
endmodule
