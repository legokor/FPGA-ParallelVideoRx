`timescale 1ns / 1ps

module dvp_receiver (
    input pclk,
    input [7:0] din,
    input href,
    input vsync,

    (* X_INTERFACE_PARAMETER = "CLK_DOMAIN pclk" *)
    (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 M_AXIS TDATA" *)
    output [7:0] tdata,
    (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 M_AXIS TLAST" *)
    output tlast,
    (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 M_AXIS TVALID" *)
    output tvalid,
    (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 M_AXIS TUSER" *)
    output tuser
);

/*
 * Rename clock
 */
wire clk;
assign clk = pclk;

/*
 * Store incoming data
 */
reg [7:0] dreg;

always @(posedge clk)
    if (href)
        dreg <= din;

reg dreg_valid;
always @(posedge clk)
    dreg_valid <= href;

/*
 * Start-of-Frame is active until the first byte after a VSYNC pulse
 */
reg sof;
always @(posedge clk)
    if (vsync)
        sof <= 1'b1;
    else if (dreg_valid)
        sof <= 1'b0;


/*
 * Set stream outputs
 */
assign tdata = dreg;
assign tlast = dreg_valid & ~href;             // Activate TLAST when HREF ends
assign tvalid = dreg_valid;
assign tuser = sof & dreg_valid;               // Activate SOF only for a single transaction

endmodule
